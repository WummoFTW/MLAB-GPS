module CA_master(
    input               rst,
    input         [4:0] prn_select,

    output reg [1022:0] CA_code 

);

always_comb begin
        case (prn_select)
            6'd1: CA_code = 1023'b110010000011100101001001111001010001001111101010110100010001010101011001000111101001111110110111001101111100101010100001000000001110101001000100110111100000111101011100110011110110000000101111001111101010011000101101110001101111010100010101100000100000000100000011000111011000000111000110111111111010011101001011011000010101011000100111001011011101100011101110111100001101100001100100100100000110110100101101111000101110000001010010011111100000101010111001111101011111001100110001110001101101010101101100011011101110000000000010110011011001110110100000101010111010111010010100011100111000100101000101001011010000101011011010110110001110011110110010000111111001011010001000011111010101110011001001001001011111111110000111110111100011011100101100001110010101000010100101011111100011110110100111011001111110111110100011000111110000000100101000101101000100010011011000000111011010001101000100100011100010110011001001111001101111110011001010011010011010111100110110101001110111100011010100010000100010010011100001110010100010000;  // PRN1 taps
            6'd2: CA_code = 1023'b111001000011100000111110100110010110111111001011001011111111010010110000100010001011000111100011000001100111000010001110001000111010011110000010110100001101001011110000111000001111100011011100110001101011100000001111000110100010111001000110011001101101001100000101111000100100101010001100000010101010000010011110000010010111111111111011101010110101010000010101001010101010000100100011001000010100001001010011011100000011100101010100110111000001111011101100000010001000101101011100110101001001100100111011011111010110000010010111100111000010110000110100011010110000001001011101100010100101101110100101101100111110000010001000101011010010100011101001110110010010001111101011111011110110001110101110101001101111001101010010111010111100000111101111101101111010001111100110110111100010000101101011010000111100110010110011000001100001000011111101011001111101001100111010100010111101000011001111101000001001111010011001011111011100101101101001111011001110011110010110111001100110101111101111011010010100101101000000101000011001000;  // PRN2 taps
            6'd3: CA_code = 1023'b111100100011100010000101001001110101000111011011110100001000010001000100010000111010011011001001000111101010110110011001101100100000000101100001110101111011110000100110111101110011010010100101001110101011011100011110011101000100001111101111100101001011101000000110100111011010111100101001011100000010001101110100101111010110101100010101111010000001001001101000110001111001110110000000111110011101010111101100001110010101010111010111100011010001010011000110111101100011011101101010010111011011111100010000111101001010000011011101001101001111010011111110000010110101010000111001011101101011001011010101111111001001010110100001100101111100111101000100001110100111100101011010001001100111110000011101011001110111010100111000011100010011101010001110011100001101101001000111000011100010111100001101010100011101110100111011000010101001100000010111100011100001100011001011110000001110100100001010001101111100011110110001001100000101000010111000001011100100001111000110110001101110001001110010111111001111110010010000000101000100100;
            6'd4: CA_code = 1023'b111110010011100011011000111110000100111011010011101011110011110000111110001001100010110101011100000100101100001100010010011110101101001000010000010101000000101101001101111111001101001010011001110001001011000010010110110000110111010100111011011011011000111010000111001000100101110111111011110011010110001010000001111001110110000101100010110010011011000101010110001100010000001111010001000101011001111000110011100111011110001110010110001001011001000111010011100010010110100101110001000110010010110000000101001100000100000011111000011000001001100010011011001110110111111100001011000010001100011001101101110110110010111100110101000010101011110010010010110010111101010000000010110000101111001111000100100001111011011000001101001111000100011100111110100100110110011010010111111001100010100000111110010110001101010111111111000011001101110001100010111110101111110100110011011001010111010111101000111111000110101100100101000101101001110101010000110011110001000111101110110101101010011010111100001101100010011101111000010011101010010;
            6'd5: CA_code = 1023'b100101101100010001101100010101110001111010101110111110011011111010100011111011100100010110010011101011110110010010000110000000011100000011100111101111010010011011011101100101101111001111011100100110110110011100010000000100100101000111111110000111001011011010001110011101110100011011100010100000010110100001001101011110001111110001001100110000000101111111110011000101100101111100100100101010011111010101100101101001001100000001100000010111011010000100011110110110100011011000011101001000011100001100110001000010100100000100110100101000101101101010101010001110101110111000010110010101011111111100010011111100100100100000001101101110000101011110110111110000100110011101111000111110101010011101001110100000111010011100111110100011101111000111000100100001011101110110010010011001100000011011010001110101110101000111000000110100001110000101010000001111110011011110110101010100100011000000001100100101011101001111100100110011010010100011010101001111000000111110010001110101010110001011100111101011010100110100000100110101001110010;
            6'd6: CA_code = 1023'b110010110100011010101100010000000110100101101001001110111010000101001101111100001101110011110001010010100010011110011101101000110011001011010011011000010100011000110000010011000011000100100101000101000101100010010001111100000111110000110011101010011000100011000011010101110010100100011110001101011100011100011101000001011010101011001110010111011001011110011011110110011110001010000011001111011000111001110111010100110010100101001101110011011100101100111111100111110110100111001010101001110001001000010101110011110011000000001100101010111000111110110001001000111010001000011100100110010110000010001110110111000100000111100011000111010111000011101011001101111101101100010011101011001001111001101101011101011101111100001110010000111010001010011011111010011110010101111101010100100011110011010000000110111001001110000010111000011110000011000001001000100110101010001100001011000001100101101011101011010110000100001111111010000010000101100110010001100011011111000101010111110110011011110110100111101111111110110010001011101111001;
            6'd7: CA_code = 1023'b100101100111111111010010011010010000111001010001100010010100101001101000111110010110111110001011011100100111001100010111101001110010001111100000110100111111000011001010010110101000101000100000100101000111011001111110011111111111100000001100011101011011010111110001100100101110001110011000000000101000001011111001011011000001001000001111100001100010001000011110001010101111110011111100001111100100101000101100110010000100001100110001010101111000101111100000011001100000000010010100000001111110100010111000110010100000101110011100011110100001000011001010011011001000101011101010101111001000111101011100100001110110000100110111010111111111101001010100100110001101011010110001111001010001010010001111000001011100110110100100011101011001000000000011111111000111110001000010011010000110000011000011110001101101100111001100010110000000101110111001111101001100011011111110011010111111010110011011110011001111101110101001010101101111100100010111100110000101111110110001010111001111111101110010000110101001110110110001000011001100100;
            6'd8: CA_code = 1023'b110010110001101101110011010111110110000100010110100000111101101100101000011110110100100111111101001001001010110001010101011100000100001101010000110101100010110100111011101010100000110111011011000100111101000000100110110001101010100011001010100111010000100101111100101001011111101110100011011101000011001001000111000011111101110111101111111111101010100101101101010001111011001101101111011101100101000111010011111001010110100011100101010010001101111001000000110000010111001010001110001101000000011111010001001011110001010101011000110001111110101010000001000010001001000001100010111011011101100010101001011001101101010101111110011011101010011000011010100110101000001111110111001000110100011110001101101101101110101001000011001111100001001001111000010101010011010110010101010101010000111111011001000100110101011110000100101001011001010110110101110001111001001000101001101100001111101110100000000000011111010100101001001001011100100110000111000101000001111111010101000110111010100000111100010001010001011111101000110000101110010;
            6'd9: CA_code = 1023'b111001011010100100100011110001000101011010110101000001101001001110001000001110100101101011000110000011111100001111110100000110111111001100001000110101001100001111000011010100100100111000100110110100000000001100001010100110100000000010101001111010010101011100111010001111100111011110111110110011110110101000011000001111100011101000011111110000101110110011010100111100010001010010100110110100100101110000101100011100111111110100001111010001110111010010010000100100101100101110000011001011011111000001100101110111011001101000111010100110010001011110100100101110101001110100100110110001010111001101010011100101100000111101011010111101100000100000111101100110111010100101010100010000000110111000001100111011110111100110110000100110111101001101000101100000011001000101111110110010111011100001010100011110011001000010100000110110110101101010110011110111100011100001000010010111010111110010111101111001110111001001101001000111000101000111001111010100100011111111100111001110000000001110011011011010101101001011000100001001011111001;
            6'd10: CA_code = 1023'b110100010010100010011100001101101000010000001000010001110110011011010010001100000010110111100111101011001111110100000010100001011010001011100100100111110001110001100111111001000000111110001110010101010001011001110101110001000001101111101101011110100100001011111110110111100101001011101010101000110000111100101000000101010000100001100001101101100101010011110011010010111000000000111011101000011000101011011101110111101010010111101011110010001010110101110000010100011111111011001110010100000100000010000110011000010100101011010010100111100010010010101101101100100101100100100000100000010000011000100111011100111111011111111111011010101110101011110110001101110011110101110010100011011000011011101101101111010101000110100000110111110001110110001111010110100111100100100100001001111010111001010100110000100010111010011110110010111010010111000011001010101111001101010101011101110110010001100000111100001110001111001111111111110101011010100001100001000010100000101011010000011111111110010100011110111011110010101001100011000000000;
            // Add cases for other PRN numbers (up to PRN 32)
            default: CA_code = 1023'b110010000011100101001001111001010001001111101010110100010001010101011001000111101001111110110111001101111100101010100001000000001110101001000100110111100000111101011100110011110110000000101111001111101010011000101101110001101111010100010101100000100000000100000011000111011000000111000110111111111010011101001011011000010101011000100111001011011101100011101110111100001101100001100100100100000110110100101101111000101110000001010010011111100000101010111001111101011111001100110001110001101101010101101100011011101110000000000010110011011001110110100000101010111010111010010100011100111000100101000101001011010000101011011010110110001110011110110010000111111001011010001000011111010101110011001001001001011111111110000111110111100011011100101100001110010101000010100101011111100011110110100111011001111110111110100011000111110000000100101000101101000100010011011000000111011010001101000100100011100010110011001001111001101111110011001010011010011010111100110110101001110111100011010100010000100010010011100001110010100010000; // Default to PRN1 taps
        endcase
    end

endmodule